
package shift_reg_config;
    import  uvm_pkg ::*;
`include "uvm_macros.svh";

    class shift_reg_config_class extends uvm_object;
    `uvm_object_utils(shift_reg_config_class);

    function new (string name = "shift_reg_config_class");
    super.new(name);
    endfunction
    endclass
    
endpackage : shift_reg_config

